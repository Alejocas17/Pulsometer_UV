** Profile: "SCHEMATIC1-alejocas"  [ C:\Users\alejo\Desktop\Universidad Del Valle\Sexto Semestre\Circuitos Electronicos\OrCad\filtro-pspicefiles\schematic1\alejocas.sim ] 

** Creating circuit file "alejocas.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.3\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 15s 0 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
